library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity memory is
    generic (
        node_address_size   : natural;
        node_size           : natural;
        nodes_to_write      : natural;
        nodes_in_parallel   : natural
    );
    port(
        clk, write_in           : in  std_logic; 
        node_data_write         : in  std_logic_vector(nodes_to_write * node_size - 1 downto 0); 
        node_addresses_write    : in  std_logic_vector(node_address_size - 1 downto 0);
        node_addresses_read     : in  std_logic_vector(nodes_in_parallel * node_address_size - 1 downto 0);
        node_data_read          : out std_logic_vector(nodes_in_parallel * node_size - 1 downto 0)
    ); 
end memory;

architecture arch of memory is

type ram_array is array (0 to (2**node_address_size) - 2) of std_logic_vector (node_size - 1 downto 0);

signal ram_data: ram_array :=(
    b"0010000000010000000",
    b"0110001110110000000",
    b"0100001111010000000",
    b"0011110100110000000",
    b"0101101001110000000",
    b"0111001111100000000",
    b"0110111010110000000",
    b"0101001100110000000",
    b"0100011010110000000",
    b"0001000000110000000",
    b"0110001111011101110",
    b"0110010011110000000",
    b"0000101111010000000",
    b"0000000000110000000",
    b"1000000000000000001",
    b"0111011010110000000",
    b"0100000111010000000",
    b"0001000000110000000",
    b"0011111000110000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"0110001111001101110",
    b"0100101101010000000",
    b"1000000000000000010",
    b"0001100001010000000",
    b"0101001000110000000",
    b"0000110000010000000",
    b"0101101111010000000",
    b"0100010101110000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"0000101001010000000",
    b"0001100001000000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"0101000101110000000",
    b"0000101001010000000",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0101101101110000000",
    b"0000101100011111000",
    b"0001100000010000000",
    b"0000101010000000000",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"0000101011110000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"0111011000110000000",
    b"0110110001010000000",
    b"0101001001110000000",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"0111010000110000000",
    b"0110001001010000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0001100000110000000",
    b"0101001101110000000",
    b"0100101000110000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0100101010100000000",
    b"0101001011100000000",
    b"1000000000000000011",
    b"1000000000000000000",
    b"0101001000110000000",
    b"1000000000000000001",
    b"0000000000110000000",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0100100110110000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"0100011011010000000",
    b"1000000000000000010",
    b"0110011001000000000",
    b"0000101001010000000",
    b"0000101011110000000",
    b"0111010010110000000",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"0001100000110000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"0100010110100000000",
    b"0110111011110000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0100100101010000000",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000000",
    b"1000000000000000000",
    b"0100001011100000000",
    b"0011111011110000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"0001100000110000000",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0110010000100000000",
    b"0101001011110000000",
    b"1000000000000000010",
    b"0110111010000000000",
    b"0100100110110000000",
    b"1000000000000000001",
    b"0011101110110000000",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"0110111010110000000",
    b"1000000000000000001",
    b"0101110100000000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0001100001000000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"0110101101100000000",
    b"0111010110010000000",
    b"0001000000110000000",
    b"0110010010010000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"0110110100100000000",
    b"0100010001010000000",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0011101110110000000",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0101101111110000000",
    b"0010100000010000000",
    b"1000000000000000001",
    b"0101110000010000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000001",
    b"0100100110110000000",
    b"0100011000110000000",
    b"0110110010110000000",
    b"0100001010010000000",
    b"0111001011110000000",
    b"1000000000000000001",
    b"0001100001000000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"0111010001000000000",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0000101110110000000",
    b"0111001101110000000",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"0100001101010000000",
    b"0000101110110000000",
    b"1000000000000000010",
    b"0101110000010000000",
    b"0100000111010000000",
    b"1000000000000000001",
    b"0111001011010000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"0100101001110000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0011110100110000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"0101101101110000000",
    b"0110010010100000000",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"0011000000110000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"0101000111010000000",
    b"1000000000000000001",
    b"0110010101110000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000011",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000000",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000010",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001",
    b"1000000000000000001"
);

begin

    process(clk, write_in)
    begin
        if rising_edge(clk) and write_in = '1' then 
            Data_serialize : for i in 0 to nodes_to_write - 1 loop
                ram_data(to_integer((i * node_address_size) + unsigned(node_addresses_write(node_address_size - 1 downto 0)))) 
                        <= 
                        node_data_write(node_size * (i + 1) - 1 downto node_size * i);
            end loop Data_serialize;
        end if;
    end process;

    Data_fetch : for i in 0 to nodes_in_parallel - 1 generate

    constant node_data_end        : natural := node_size * (i + 1) - 1;
    constant node_data_start      : natural := node_size * i;
    constant node_address_end        : natural := node_address_size * (i + 1) - 1;
    constant node_address_start      : natural := node_address_size * i;

    begin
        node_data_read(node_data_end downto node_data_start) <= ram_data(to_integer(unsigned(node_addresses_read(node_address_end downto node_address_start))));
    end generate Data_fetch;

end arch;
