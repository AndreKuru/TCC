library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity register_bank is
    generic (
        node_address_size   : natural;
        node_size           : natural;
        nodes_to_write      : natural;
        nodes_in_parallel   : natural
    );
    port(
        clk, write_in           : in  std_logic; 
        node_data_write         : in  std_logic_vector(nodes_to_write * node_size - 1 downto 0); 
        node_addresses_write    : in  std_logic_vector(node_address_size - 1 downto 0);
        node_addresses_read     : in  std_logic_vector(nodes_in_parallel * node_address_size - 1 downto 0);
        node_data_read          : out std_logic_vector(nodes_in_parallel * node_size - 1 downto 0)
    ); 
end register_bank;

architecture arch of register_bank is

type ram_array is array (0 to (2**node_address_size) - 2) of std_logic_vector (node_size - 1 downto 0);

signal ram_data: ram_array :=(
    b"001000000001000000000",
    b"010100100111000101000",
    b"010000111101000000000",
    b"010100100110000101000",
    b"011101000010000000000",
    b"011100111110000000000",
    b"011011101011000000000",
    b"011000111011000000000",
    b"000010110001111100011",
    b"011001101111000000000",
    b"000100000001000000000",
    b"011001001111000000000",
    b"000010111101000000000",
    b"000000000001000000000",
    b"100000000000000000000",
    b"010100011011000000000",
    b"010110100111000000000",
    b"100000000000000000000",
    b"011101010111010111100",
    b"001111001111000000000",
    b"100000000000000000001",
    b"010000100111000000000",
    b"000110000011000000000",
    b"100000000000000000001",
    b"000010100101000000000",
    b"010100100011000000000",
    b"000011000001000000000",
    b"010001010111000000000",
    b"010010011101000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010111000000101011000",
    b"100000000000000000000",
    b"000100000001000000000",
    b"010111010110000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010001001000000000000",
    b"100000000000000000010",
    b"100000000000000000000",
    b"001111010110000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010000100001000000000",
    b"000011000011000000000",
    b"100000000000000000000",
    b"001111101111000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"011011011111000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"010100100111000000000",
    b"100000000000000000001",
    b"011011001010000000000",
    b"010010110001000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011101011000010111100",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"011000111100110111010",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010010010101000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010000011011000000000",
    b"001111100011000000000",
    b"100000000000000000000",
    b"011101101101000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"001111010001000000000",
    b"010100110010000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"001111001010000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010010011011000000000",
    b"011101001011000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"011101100101000000000",
    b"011001011101000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011101011001010111100",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010110110111000000000",
    b"010100100011000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"001111100100000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011101101000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010010100001000000000",
    b"011010111111000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"011101000011000000000",
    b"010001010101000000000",
    b"000010101101000000000",
    b"010111000001000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"011101100011000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"011011100001000000000",
    b"010000101110000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011011100000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011100111111000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"000010101111000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"010111010000000000000",
    b"011101100111000000000",
    b"010001011010000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"000010110011000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"011101100011000000000",
    b"011010110110000000000",
    b"011101011001000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010100101010000101000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010001010001000000000",
    b"100000000000000000000",
    b"011011000101000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"011011000110000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"001010000001000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010110110101000000000",
    b"010001100011000000000",
    b"011011001011000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010001010101000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011001001001000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000010",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000"
);

begin

    process(clk, write_in)
    begin
        if rising_edge(clk) and write_in = '1' then 
            Data_serialize : for i in 0 to nodes_to_write - 1 loop
                ram_data(to_integer((i * node_address_size) + unsigned(node_addresses_write(node_address_size - 1 downto 0)))) 
                        <= 
                        node_data_write(node_size * (i + 1) - 1 downto node_size * i);
            end loop Data_serialize;
        end if;
    end process;

    Data_fetch : for i in 0 to nodes_in_parallel - 1 generate

    constant node_data_end        : natural := node_size * (i + 1) - 1;
    constant node_data_start      : natural := node_size * i;
    constant node_address_end        : natural := node_address_size * (i + 1) - 1;
    constant node_address_start      : natural := node_address_size * i;

    begin
        node_data_read(node_data_end downto node_data_start) <= ram_data(to_integer(unsigned(node_addresses_read(node_address_end downto node_address_start))));
    end generate Data_fetch;

end arch;
