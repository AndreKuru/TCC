library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity memory is
    generic (node_address_size  :natural;
            node_size           :natural;
            nodes_in_parallel   :natural := 3);
    port(
        clk, write_in   : in  std_logic; 
        node_addresses  : in  std_logic_vector(nodes_in_parallel * node_address_size - 1 downto 0);
        node_data_in    : in  std_logic_vector(nodes_in_parallel * node_size - 1 downto 0); 
        node_data_out   : out std_logic_vector(nodes_in_parallel * node_size - 1 downto 0)
    ); 
end memory;

architecture arch of memory is

type ram_array is array (0 to (2 ** node_address_size) - 1) of std_logic_vector (node_size - 1 downto 0);

signal ram_data: ram_array :=(
    b"1000000000000011000000010111100110000000000000000",
    b"1000000000000010110000000000000100001110101110000",
    b"1000000000000001100000000000000100010101000111101",
    b"1000000000000010100000000000000001110111101011100",
    b"1000000000000001100000000000000001100101110000101",
    b"1000000000000000010000000000000100001010111000010",
    b"1000000000000010010000000000000110110111101011100",
    b"1000000000000001100000000000000011001010001111010",
    b"1000000000000010010000000000001011101000010100011",
    b"1100000000000000000000000000000000000000000000000",
    b"1000000000000000000000000000011010010110011001100",
    b"1100000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"1000000000000010010000000000001000000111101011100",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"1100000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000",
    b"0000000000000000000000000000000000000000000000000"
);

begin

    process(clk)
    begin
        if rising_edge(clk) and write_in = '1' then 
            Data_serialize : for i in 0 to nodes_in_parallel loop
                ram_data(to_integer(unsigned(node_addresses))) <= node_data_in(
                                                                    node_size * i 
                                                                    downto 
                                                                    node_size * (i + 1) - 1);
            end loop Data_serialize;
        end if;
    end process;

    Data_fetch : for i in 0 to nodes_in_parallel generate

    signal node_data_start      : natural := node_size * i;
    signal node_data_end        : natural := node_size * (i + 1) - 1;

    begin
        node_data_out(node_data_end downto node_data_start) <= ram_data(to_integer(unsigned(node_addresses)));
    end generate Data_fetch;

end arch;