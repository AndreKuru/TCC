library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity register_bank is
    generic (
        node_address_size   : natural;
        node_size           : natural;
        nodes_to_write      : natural;
        nodes_in_parallel   : natural
    );
    port(
        clk, write_in           : in  std_logic; 
        node_data_write         : in  std_logic_vector(nodes_to_write * node_size - 1 downto 0); 
        base_address_to_write    : in  std_logic_vector(node_address_size - 1 downto 0);
        node_addresses_read     : in  std_logic_vector(nodes_in_parallel * node_address_size - 1 downto 0);
        node_data_read          : out std_logic_vector(nodes_in_parallel * node_size - 1 downto 0)
    ); 
end register_bank;

architecture arch of register_bank is

type ram_array is array (0 to (2**node_address_size) - 2) of std_logic_vector (node_size - 1 downto 0);

signal ram_data: ram_array :=(
    b"001000000001000000000",
    b"010100100011000000000",
    b"010000111101000000000",
    b"011000111011000000000",
    b"010010110101000000000",
    b"011100111110000000000",
    b"011011101011000000000",
    b"010001101011000000000",
    b"010110100111000000000",
    b"010111001011000000000",
    b"011001101000000000000",
    b"011001001111000000000",
    b"000010111101000000000",
    b"000000000001000000000",
    b"100000000000000000000",
    b"000110000001000000000",
    b"011011101010000000000",
    b"000100000001000000000",
    b"010000101110000000000",
    b"010110111011000000000",
    b"000100000001000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"000110000011000000000",
    b"010100100011000000000",
    b"000011000001000000000",
    b"010001010111000000000",
    b"010110111101000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011011011011000000000",
    b"010001011011000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"010000100101000000000",
    b"011101010001000000000",
    b"000010101100000000000",
    b"100000000000000000000",
    b"010000101001000000000",
    b"011101000011000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"011011011111000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"010100100111000000000",
    b"100000000000000000001",
    b"011101100011000000000",
    b"011011000101000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011000100110000000000",
    b"010010100011000000000",
    b"100000000000000000000",
    b"010100011001000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"011101100011000000000",
    b"010001100010000000000",
    b"011011001011000000000",
    b"000010101001000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010000011011000000000",
    b"001111101111000000000",
    b"001111001100000000000",
    b"000110000011000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"000110000001000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010010011011000000000",
    b"000100000001000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010001101101000000000",
    b"100000000000000000001",
    b"011001100100000000000",
    b"000010100101000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"010110101101000000000",
    b"100000000000000000000",
    b"011000101011000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010010010111000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011001001101000000000",
    b"011001000101000000000",
    b"010111001101000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"000000000001000000000",
    b"100000000000000000000",
    b"010001000100000000000",
    b"100000000000000000000",
    b"001111010110000000000",
    b"100000000000000000000",
    b"010010010110000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010010100001000000000",
    b"001111011001000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010100010111000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"011001000010000000000",
    b"010111011011000000000",
    b"100000000000000000001",
    b"011011101000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010001011001000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"000010100111000000000",
    b"010010011001000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010010100111000000000",
    b"010111001101000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"000010111101000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011100111111000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"000110000001000000000",
    b"001110101100000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010000111111000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010110111111000000000",
    b"010100110001000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011001010000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"001111010010000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"010110101100000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"010100100011000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"011011011100111010111",
    b"011100110111000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"011001001101000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"000110000010000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000001",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000",
    b"100000000000000000000"
);

begin

    process(clk, write_in)
    begin
        if rising_edge(clk) and write_in = '1' then 
            Data_serialize : for i in 0 to nodes_to_write - 1 loop
                ram_data(to_integer((i * node_address_size) + unsigned(base_address_to_write(node_address_size - 1 downto 0)))) 
                        <= 
                        node_data_write(node_size * (i + 1) - 1 downto node_size * i);
            end loop Data_serialize;
        end if;
    end process;

    Data_fetch : for i in 0 to nodes_in_parallel - 1 generate

    constant node_data_end        : natural := node_size * (i + 1) - 1;
    constant node_data_start      : natural := node_size * i;
    constant node_address_end        : natural := node_address_size * (i + 1) - 1;
    constant node_address_start      : natural := node_address_size * i;

    begin
        node_data_read(node_data_end downto node_data_start) <= ram_data(to_integer(unsigned(node_addresses_read(node_address_end downto node_address_start))));
    end generate Data_fetch;

end arch;
